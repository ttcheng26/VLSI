library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity counter is
port(
	  add_A: in std_logic_vector(7 downto 0);
	  add_B: in std_logic_vector(7 downto 0);
	  sum : out std_logic_vector(7 downto 0));
end counter;

architecture behavior of counter is
begin
	process(add_A)
		begin
			sum <= add_A + add_B;
	end process;
end behavior;
